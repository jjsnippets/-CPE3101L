// CPE 3101L - INTRODUCTION TO HDL
// Group 1		F 7:30 - 10:30 AM LB285TC
// LabExercise #4
// Sarcol, Joshua S.		BS CpE - 3		2025/09/19

// 
// Testbench file for mux_4_to_1_nb.v (unit test)
// 
`timescale 1 ns / 1 ps
module tb_mux_4_to_1_nb ();
